`define LENGTH 4
